



module cache
(
    WB4.master master_bus,
    WB4.slave slave_bus
);









endmodule