

module vga_controller
(
    WB4 wb.slave wb   
);




endmodule