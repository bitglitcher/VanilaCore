
interface SPI;
    logic MISO;
    logic MOSI;
    logic SCLK;
    logic [3:0] CS;
endinterface //SPI