
interface SPI;
    logic MISO;
    logic MOSI;
    logic SCLK;
endinterface //SPI