
`ifndef __DEBUG__PORT__SV__
`define __DEBUG__PORT__SV__

`define DEBUG_PORT
`define MEMORY_DEBUG_MSGS

`endif