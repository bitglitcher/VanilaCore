


ram_wb MEMORY_INST();
ram_wb MEMORY_DATA();