

//This is the implementation for the CSR Cycle counter

module csr_timer();













