
`define DEBUG_PORT