


module spi
(
    WB4.slave wb
);

//0x0000 DATA
//










endmodule