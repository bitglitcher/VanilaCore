





module feedback_latched();

logic cyc1;
logic cyc2;


logic cyc1_out;
logic cyc2_out;


initial begin
    cyc1 = 0;
    cyc2 = 0;
    cyc1_out = 0;
    cyc2_out = 0;
end



always @() begin
    
end