
module performance_counter
(
    input logic [11:0] addr,
    input logic wr,
    input  logic [31:0] din,
    output logic [31:0] dout
);















endmodule