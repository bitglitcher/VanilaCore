interface csr_int;
    
endinterface //csr_int